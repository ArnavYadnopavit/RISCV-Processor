module instruction_memory (
        input  wire         clk,
    	input  wire [9:0] pc,         
    	output reg [31:0] instruction
);
    	(* ram_style = "block" *)reg [7:0] memory [0:1023];       //1024 x 8-bit = 1 KB instruction_memory
        
    	always @(posedge clk) begin
        	instruction <= { memory[pc], memory[pc+1], memory[pc+2], memory[pc+3] };  
    	end

    	// preload program from file
    	initial begin
        	$readmemh("program.hex", memory);
    	end
endmodule

