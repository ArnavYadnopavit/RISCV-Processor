module ALU(
    input a[63:0],
    input b[63:0],
    input control[]
    output out[63:0],
    output flagzero;
)

always @(*) begin
    
end

endmodule