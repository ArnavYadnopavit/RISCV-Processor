`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 15.11.2025 18:40:29
// Design Name: 
// Module Name: dmemstaller
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module dmemstaller(
    input clk,
    input reset,
    input MemWrite,
    input MemRead,
    output reg MemStall
    );
    wire isMem;
    assign isMem=MemWrite||MemRead;
    always@(negedge clk or posedge reset or posedge isMem)begin
        if(reset)MemStall<=1'b0;
        casez(MemStall)
            1'b0:if(isMem)begin
                MemStall<=1'b1;
                end
                else MemStall<=1'b0;
            1'b1:MemStall<=1'b0;
            default:MemStall<=1'b0;        
        endcase
    end 
endmodule
