module mem_wb_reg(
        input wire clk,
        input wire reset,
		input wire [63:0] mem_data_in,     
        input wire [63:0] alu_result_in,   
        input wire [63:0] pc_in,
		input wire [4:0] rd_in,       
        input wire RegWrite_in,
        input wire MemtoReg_in,
        input wire Jump_in,
		input wire StallW,
		output reg [63:0] mem_data_out,
        output reg [63:0] alu_result_out,
        output reg [63:0] pc_out,
        output reg [4:0] rd_out,
        output reg RegWrite_out,
        output reg MemtoReg_out,
        output reg Jump_out
        

);

        always @(posedge clk or posedge reset) begin
                if (reset) begin
                        mem_data_out <= 64'b0;
                        alu_result_out <= 64'b0;
                        pc_out <= 64'b0;
                        rd_out <= 5'b0;
                        RegWrite_out <= 1'b0;
                        MemtoReg_out <= 1'b0;
                        Jump_out <= 0;
                end 
                
 			else if (StallW) begin
    				mem_data_out   <= mem_data_out;
    				alu_result_out <= alu_result_out;
    				pc_out <= pc_out;
    				rd_out <= rd_out;
    				RegWrite_out <= RegWrite_out;
    				MemtoReg_out <= MemtoReg_out;
    				Jump_out <= Jump_out;
			end

    		else begin
        			mem_data_out   <= mem_data_in;
        			alu_result_out <= alu_result_in;
        			pc_out         <= pc_in;
        			rd_out         <= rd_in;
        			RegWrite_out   <= RegWrite_in;
        			MemtoReg_out   <= MemtoReg_in;
        			Jump_out       <= Jump_in;
    		end
			
		end
	
endmodule

