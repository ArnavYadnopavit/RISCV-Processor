module pipelined_datapath(
        input  wire clk,
        input  wire reset,
        output wire [63:0] debug_pc,
        //output wire [63:0] debug_alu_result,
        //output wire [63:0] debug_alu_input1,
     //   output wire [63:0] debug_alu_input2,
     //   output wire [63:0] debug_regfile_out2,
     //   output wire [63:0] debug_imm_out,
        output wire [31:0] inst_debug
     //   output wire valid_alu_debug,
      //  output wire [4:0] debug_alu_control
);

//DECLARING WIRES
        wire [63:0] pc_out;
        wire [63:0] pc_next;

        wire [31:0] instruction;

  	wire [2:0] ALUOp;
  	wire RegWrite, ALUSrc, MemtoReg, Branch, Jump, MemRead, MemWrite;
  	wire InstType;

        wire [63:0] read_data1;
        wire [63:0] read_data2;
        wire [63:0] write_data;

        wire [63:0] imm;

        wire [63:0] alu_result;
        wire [4:0]  ALUControlPort;
        wire branch_D;
        wire valid;

        wire [63:0] mem_data;
        
        //wire take_branch;
        
        wire [63:0] if_id_pc_out;
	wire [31:0] if_id_instruction_out;
	
  	wire [6:0] opcode = if_id_instruction_out[6:0];
  	wire [4:0] rd = if_id_instruction_out[11:7];
  	wire [2:0] func3 = if_id_instruction_out[14:12];
  	wire [4:0] rs1 = if_id_instruction_out[19:15];
  	wire [4:0] rs2 = if_id_instruction_out[24:20];
  	wire [6:0] func7 = if_id_instruction_out[31:25];
  	wire op5 = opcode[5];
  	wire func75 = func7[5];
  	wire func70 = func7[0];
  	
  	wire [63:0] id_ex_pc_out, id_ex_rs1_out, id_ex_rs2_out, id_ex_imm_out;
  	wire [4:0] id_ex_rd_out;
  	wire [2:0] id_ex_func3_out, id_ex_ALUop_out;
  	wire [6:0] id_ex_opcode_out;
  	wire id_ex_func75_out,id_ex_func70_out, id_ex_op5_out;
 	wire id_ex_ALUSrc_out, id_ex_RegWrite_out, id_ex_MemtoReg_out;
  	wire id_ex_Branch_out, id_ex_Jump_out, id_ex_MemRead_out, id_ex_MemWrite_out, id_ex_InstType_out;
  	wire [4:0] id_ex_rs1_E_out;
	wire [4:0] id_ex_rs2_E_out;
	wire DivStalled;
	wire MemStall;
	wire Divreset;
	
	
	wire [63:0] ex_mem_pc_out, ex_mem_alu_result_out, ex_mem_rs2_out;
	wire [2:0]  ex_mem_func3_out;
  	wire [4:0] ex_mem_rd_out;
 	//wire ex_mem_branchAlu_out;
 	wire ex_mem_RegWrite_out, ex_mem_MemRead_out, ex_mem_MemWrite_out;
  	wire ex_mem_MemtoReg_out, ex_mem_Jump_out;
  	//wire  ex_mem_Branch_out;
  	
  	wire [63:0] mem_wb_mem_data_out, mem_wb_alu_result_out, mem_wb_pc_out;
  	wire [4:0] mem_wb_rd_out;
  	wire mem_wb_RegWrite_out, mem_wb_MemtoReg_out,mem_wb_Jump_out;
  	
	wire [63:0] branchpc;
	
	wire StallD, StallF,StallE,StallM,FlushD, FlushE;
 	wire [1:0] ForwardAE, ForwardBE;
 	wire [63:0] BranchD_in1,BranchD_in2;
 	wire [1:0] BranchForwardAE,BranchForwardBE;
 	
 	wire [63:0] srcA_E, srcB_E_pre, srcB_E;
 	
 	wire PcSrc;
	assign PcSrc = Jump || (Branch && branch_D);
	
	assign FlushD = PcSrc;



	
        //instruction_memory IM (
          //      .clk(clk),
           //     .pc(pc_out),
           //     .instruction(instruction)
        //);
        
	program_counter PC (
  		.clk(clk),
  		.reset(reset),
  		.stall(StallF),
  		.pc_next(pc_next),
  		.pc_out(pc_out)
	);
          
    	imem_ip IM(
        	.clka(~clk),
        	.ena(1'b1),
        	.wea(4'b0),
        	.addra(pc_out[15:2]),
        	.dina(32'd0),
        	.douta(instruction)
    	);
        
	if_id_reg IF_ID (
  		.clk(clk),
  		.reset(reset),
  		.enable(~StallD),
  		.FlushD(FlushD),
  		.instruction_in(instruction),
  		.pc_in(pc_out),
  		.instruction_out(if_id_instruction_out),
  		.pc_out(if_id_pc_out)
	);

	ControlUnit CU (
        	.opcode(opcode),
        	.func3(func3),   
        	.ALUOp(ALUOp),
        	.RegWrite(RegWrite),
        	.ALUSrc(ALUSrc),
        	.MemRead(MemRead),
        	.MemWrite(MemWrite),
        	.MemtoReg(MemtoReg),
        	.Branch(Branch),
        	.Jump(Jump),
        	.InstType(InstType)
	);


        ImmGen IG (
                .inst(if_id_instruction_out),
                .imm(imm)
        );

        reg_file RF (
                .clk(~clk),
                .reset(reset),
                .reg_write(mem_wb_RegWrite_out),
                .rs1(rs1),
                .rs2(rs2),
                .rd(mem_wb_rd_out),
                .write_data(write_data),
                .read_data1(read_data1),
                .read_data2(read_data2)
        );
        //New muxes added for branch comparing regs forwarding
        mux3 BranchD_A (
            .a(read_data1),
            .b(alu_result),
            .c(write_data),
            .sel(BranchForwardAE),
            .y(BranchD_in1)
        );
        
        mux3 BranchD_B (
            .a(read_data2),
            .b(alu_result),
            .c(write_data),
            .sel(BranchForwardBE),
            .y(BranchD_in2)
        );
        
        
        
	Branch_D brD (
  		.rs1D_data(BranchD_in1),
  		.rs2D_data(BranchD_in2),
  		.pc(if_id_pc_out),
  		.imm(imm),
  		.func3(func3),
  		.branch_dec(branch_D),
  		.branchpc(branchpc)
	);
        
        id_ex_reg ID_EX (
                .clk(clk),
                .reset(reset),
                .StallE(StallE),
                .FlushE(FlushE),
                .pc_in(if_id_pc_out),
                .rs1_D_in(rs1),
                .rs2_D_in(rs2),
                .rs1_data_in(read_data1),
                .rs2_data_in(read_data2),
                .imm_in(imm),
                .rd_in(rd),
                .func3_in(func3),
                .opcode_in(opcode),
                .func70_in(func70),
                .func75_in(func75),
                .ALUop_in(ALUOp),
                .op5_in(op5),
                .ALUSrc_in(ALUSrc),
                .RegWrite_in(RegWrite),
                .MemtoReg_in(MemtoReg),
                .Branch_in(Branch),
                .Jump_in(Jump),
                .MemRead_in(MemRead),
                .MemWrite_in(MemWrite),
                .InstType_in(InstType),
                .pc_out(id_ex_pc_out),
                .rs1_E_out(id_ex_rs1_E_out),
                .rs2_E_out(id_ex_rs2_E_out),
                .rs1_data_out(id_ex_rs1_out),
                .rs2_data_out(id_ex_rs2_out),
                .imm_out(id_ex_imm_out),
                .rd_out(id_ex_rd_out),
                .func3_out(id_ex_func3_out),
                .opcode_out(id_ex_opcode_out),
                .func70_out(id_ex_func70_out),
                .func75_out(id_ex_func75_out),
                .ALUop_out(id_ex_ALUop_out),
                .op5_out(id_ex_op5_out),
                .ALUSrc_out(id_ex_ALUSrc_out),
                .RegWrite_out(id_ex_RegWrite_out),
                .MemtoReg_out(id_ex_MemtoReg_out),
                .Branch_out(id_ex_Branch_out),
                .Jump_out(id_ex_Jump_out),
                .MemRead_out(id_ex_MemRead_out),
                .MemWrite_out(id_ex_MemWrite_out),
                .InstType_out(id_ex_InstType_out)
        );
        
  	ALUControl ALUC (
    		.op5(id_ex_op5_out),
    		.func70(id_ex_func70_out),
    		.func75(id_ex_func75_out),
    		.func3(id_ex_func3_out),
    		.AluOp(id_ex_ALUop_out),
    		.AluControlPort(ALUControlPort)
  	);
  	
  	//New Unit added for stalling div
  	DivStaller DIVSTALL(
  	     .clk(clk),
  	     .reset(reset),
  	     .AluControlPort(ALUControlPort),
  	     .DivStalled(DivStalled),
  	     .Divreset(Divreset)
  	);
  	
  	// muxes needed for ALU
  	
	mux3 muxA (
    		.a(id_ex_rs1_out),
    		.b(write_data),
    		.c(ex_mem_alu_result_out),
    		.sel(ForwardAE),
    		.y(srcA_E)
	);

	mux3 muxB (
	    .a(id_ex_rs2_out),
	    .b(write_data),
	    .c(ex_mem_alu_result_out),
	    .sel(ForwardBE),
	    .y(srcB_E_pre)
	);

	// ALUSrc select
	mux2 muxALUSrc (
	    .a(srcB_E_pre),
	    .b(id_ex_imm_out),
	    .sel(id_ex_ALUSrc_out),
    	    .y(srcB_E)
	);

	ALU ALU64 (
	        .clk(clk),
	        .Divreset(Divreset),
    		.a(srcA_E),
    		.b(srcB_E),
    		.control(ALUControlPort),
    		.out(alu_result),
    		.valid(valid),
    		.InstType(id_ex_InstType_out)
	);
	
	dmemstaller DMSTALL(
	   .clk(clk),
	   .reset(reset),
	   .MemWrite(ex_mem_MemWrite_out),
	   .MemRead(ex_mem_MemRead_out),
	   .MemStall(MemStall)	   
	);

  	ex_mem_reg EX_MEM (
    		.clk(clk),
    		.reset(reset),
    		.StallM(StallM),
    		.pc_in(id_ex_pc_out),
    		.func3_in(id_ex_func3_out),
    		.alu_result_in(alu_result),
    		//.branchAlu_in(branchAlu),
    		.alu_input2_in(id_ex_rs2_out),
    		.rd_in(id_ex_rd_out),
    		.RegWrite_in(id_ex_RegWrite_out),
    		.MemRead_in(id_ex_MemRead_out),
    		.MemWrite_in(id_ex_MemWrite_out),
    		.MemReg_in(id_ex_MemtoReg_out),
    		.Branch_in(id_ex_Branch_out),
    		.Jump_in(id_ex_Jump_out),
    		.pc_out(ex_mem_pc_out),
    		.func3_out(ex_mem_func3_out),
    		.alu_result_out(ex_mem_alu_result_out),
    		//.branchAlu_out(ex_mem_branchAlu_out),
    		.alu_input2_out(ex_mem_rs2_out),
    		.rd_out(ex_mem_rd_out),
    		.RegWrite_out(ex_mem_RegWrite_out),
    		.MemRead_out(ex_mem_MemRead_out),
    		.MemWrite_out(ex_mem_MemWrite_out),
    		.MemReg_out(ex_mem_MemtoReg_out),
    		//.Branch_out(ex_mem_Branch_out),
    		.Jump_out(ex_mem_Jump_out)
  	);


  	dmem_top DMEM (
    		.clk(clk),
    		.we(ex_mem_MemWrite_out),
    		.re(ex_mem_MemRead_out),
    		.data(ex_mem_rs2_out),
    		.addr(ex_mem_alu_result_out),
    		.func3(ex_mem_func3_out),
    		.out_data(mem_data)
  	);
        
  	mem_wb_reg MEM_WB (
    		.clk(clk),
    		.reset(reset),
    		.mem_data_in(mem_data),
    		.alu_result_in(ex_mem_alu_result_out),
    		.pc_in(ex_mem_pc_out),
    		.rd_in(ex_mem_rd_out),
    		.RegWrite_in(ex_mem_RegWrite_out),
    		.MemtoReg_in(ex_mem_MemtoReg_out),
    		.Jump_in(ex_mem_Jump_out),
    		.mem_data_out(mem_wb_mem_data_out),
    		.alu_result_out(mem_wb_alu_result_out),
    		.pc_out(mem_wb_pc_out),
    		.rd_out(mem_wb_rd_out),
    		.RegWrite_out(mem_wb_RegWrite_out),
    		.MemtoReg_out(mem_wb_MemtoReg_out),
    		.Jump_out(mem_wb_Jump_out)   
  	);
  	
  	wire [1:0] wb_sel;

	assign wb_sel =
		mem_wb_MemtoReg_out ? 2'b01 :   // load
		mem_wb_Jump_out     ? 2'b10 :   // JAL/JALR link address
                            	      2'b00;    // ALU result

	wire [63:0] link_val;
	assign link_val = mem_wb_pc_out + 64'd4;

  	
	mux3 wb_mux (
    		.a(mem_wb_alu_result_out),   // sel = 00
    		.b(mem_wb_mem_data_out),     // sel = 01
    		.c(link_val),                // sel = 10
    		.sel(wb_sel),
    		.y(write_data)
	);



	HazardDetection HDU (
  		.rs1_D(rs1),
  		.rs2_D(rs2),
  		.rs1_E(id_ex_rs1_E_out),
  		.rs2_E(id_ex_rs2_E_out),
  		.rd_E(id_ex_rd_out),
  		.rd_M(ex_mem_rd_out),
  		.rd_W(mem_wb_rd_out),
  		.opcode_E(id_ex_opcode_out),
  		//.PCSrc_E(1'b0), 
  		.regwrite_E(id_ex_RegWrite_out),
  		.regwrite_M(ex_mem_RegWrite_out),
  		.regwrite_W(mem_wb_RegWrite_out),
  		.MemtoregE(id_ex_MemtoReg_out),
  		.MemtoregM(ex_mem_MemtoReg_out),
  		.DivStalled(DivStalled),
  		.MemStall(MemStall),
  		.StallD(StallD),
  		//.FlushD(FlushD), 
  		.FlushE(FlushE),
  		.StallE(StallE),
  		.StallM(StallM),
  		.ForwardAE(ForwardAE),
  		.ForwardBE(ForwardBE),
  		.StallF(StallF),
  		.BranchForwardAE(BranchForwardAE),
  		.BranchForwardBE(BranchForwardBE)
);

	wire [63:0] pc_plus4;
	//wire [63:0] jal_target;
	wire [63:0] jalr_target;
	wire [1:0]  pc_sel;

	assign pc_plus4      = pc_out + 64'd4;
	//assign jal_target    = if_id_pc_out + imm;
	assign jalr_target   = read_data1 + imm + 64'd4;

	assign pc_sel[1] = Jump;
	assign pc_sel[0] = (Branch && branch_D) || (Jump && (opcode == 7'b1100111));

	mux4_64 mux_pc_next (
	    	.a(pc_plus4),
    		.b(branchpc),
    		.c(branchpc),
    		.d(jalr_target),
    		.sel(pc_sel),
    		.y(pc_next)
	);

	/*
        assign write_data = ((opcode == 7'b1101111) ||     // JAL
                     (opcode == 7'b1100111)) ? pc_out :  // JAL / JALR
                    (MemtoReg) ? mem_data :              // load
                                 alu_result;             // ALU result (includes LUI)


        

        assign take_branch = (Branch && branch_D) || Jump;
        wire [63:0]jumpimm;
        assign jumpimm=imm<<1;
        assign pc_next = take_branch ? 
                    ((Jump && (opcode == 7'b1100111)) ? (read_data1 + imm) :     // JALR
                     (Jump && (opcode == 7'b1101111)) ? (pc_out - 64'd4 + jumpimm) : // JAL
                     (pc_out - 64'd8 + jumpimm))                                     // other branch
                 : (opcode == 7'b0010111) ? imm                                       // AUIPC
                 : (pc_out + 64'd4);                                                  // normal PC increment



        
        //always @(posedge clk,posedge reset)begin
        //    if (reset) 
        //        stall<=1'b0;
        //    if(opcode== 7'b0000011 | opcode==7'b1100011 | opcode==7'b1101111 | opcode==7'b1100111)
        //        stall=~stall;
        //end
        */
        
        assign debug_pc = pc_out;
       // assign debug_alu_result = alu_result;
        assign inst_debug=instruction;
       // assign debug_alu_input1=read_data1;
       // assign debug_regfile_out2=read_data2;
      //  assign debug_imm_out=imm;
      //  assign debug_alu_input2=ALUSrc ? imm : read_data2;
      //  assign valid_alu_debug=valid;
      //  assign debug_alu_control=ALUControlPort;


endmodule

